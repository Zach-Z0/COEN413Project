/*

Wrapper class

Takes the DUT inputs/outputs delcared in "calc2_top" and equates them to interface signals

Zachary Zazzara (40096894)

Created on: March 29th, 2024
*/

module wrapper (tb_if interf);
 calc2_top DUT (
    //TODO
    //Connect DUT inputs/outputs to interface here!
    //"INTERFACE NAME" -> "DUT INTERNAL NAME"
    //The declaration from calc2_top.v is not clear. Some of the signals expected aren't in the documentation.
    // Need to email TA for help. 
 );
endmodule