/*

Monitor class for the testbench, watches the DUT outputs and passes the results up into the scoreboard/checker.
Only needs to monitor the actual OUTPUTS of the DUT.

Zachary Zazzara (40096894)
zexi si (40175054)

Created on: March 30th, 2024
*/

class moni;
    //TODO
endclass