/*

Scoreboard class, Probably will also have the checker mixed in with it? I'm not super sure yet, I need to think about how to
structure this and how I can/will need to handle mail from the agent mail arriving out of sync with the monitor mail.


zexi si (40175054 )
zachary zazzara (40096894)
*/

class tb_scb;
    //TODO
endclass: tb_scb